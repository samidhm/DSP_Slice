`timescale 1ns / 1ps

module tb_dsp6_fp32();

reg clk;
reg enable;
reg clr;
reg [3:0] funct;
reg [31:0] chainin;
reg accumulate;
reg [31:0] ax;
reg [31:0] ay;
reg [31:0] az;
wire [31:0] chainout;
wire [31:0] resulta_flopped;

dsp_slice_fp32 dsp_slice(clk, enable, clr, funct, chainin, accumulate, ax, ay, az, chainout, resulta_flopped );

initial begin
clk = 0;
repeat(40)
#10 clk = ~clk; #10 $finish;
end

initial begin
clr=1;
#5 clr=0;
end


initial begin
#30  funct= 4'b0000; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0001; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0010; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0011; accumulate = 1'b1; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0100; accumulate = 1'b1; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0101; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0110; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b0111; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b1000; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b1001; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b1010; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;
#20  funct= 4'b1010; accumulate = 1'b0; chainin = 32'b00111111010110100101011100101111 ; ax= 32'b11000000110100011100001011110010 ; ay= 32'b00111110000111111111010001001101; az= 32'b00111111010110100101011100101111;

end




endmodule
